`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:41:23 06/01/2018 
// Design Name: 
// Module Name:    car 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module car(
	// inputs 
	
	// outputs
	
    );

	reg [7:0] color;
	reg is_moving;
	reg [1:0] road_num; // starting from up is 0, clockwise
	reg [1:0] lane_num; // starting from up is 0, clockwise
	
endmodule
